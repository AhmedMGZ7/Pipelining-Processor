library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity ALU is
  port (
    clk : in std_logic
  );
end entity ALU;
architecture ALUarc of ALU is
    begin
end architecture;