library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity ForwardingUnit is
  port (
    clk : in std_logic
  );
end entity ForwardingUnit;
architecture ForwardingUnitarc of ForwardingUnit is
    begin
end architecture;