library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity load_use_detection is
  port (
    clk : in std_logic
  );
end entity load_use_detection;
architecture load_use_detectionarc of load_use_detection is
    begin
end architecture;